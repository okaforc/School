LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY mux2_32bit IS
    PORT (
        mu_In0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        mu_In1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        mu_s : IN STD_LOGIC;
        mu_Z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END mux2_32bit;

ARCHITECTURE Behavioral OF mux2_32bit IS
BEGIN
    mu_Z <= mu_In0 AFTER 2 ns WHEN mu_S = '0' ELSE
        mu_In1 AFTER 2 ns WHEN mu_S = '1'ELSE
        x"00000000";
END Behavioral;

