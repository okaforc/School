-- Michael Manzke
-- michael.manzke@cs.tcd.ie
-- 17th November 2021
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ctrl_mem IS
    PORT (
        IN_CAR : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
        FL : OUT STD_LOGIC; -- 0
        RZ : OUT STD_LOGIC; -- 1
        RN : OUT STD_LOGIC; -- 2
        RC : OUT STD_LOGIC; -- 3
        RV : OUT STD_LOGIC; -- 4
        MW : OUT STD_LOGIC; -- 5
        MM : OUT STD_LOGIC; -- 6
        RW : OUT STD_LOGIC; -- 7
        MD : OUT STD_LOGIC; -- 8
        FS : OUT STD_LOGIC_VECTOR(4 DOWNTO 0); -- 9 to 13
        MB : OUT STD_LOGIC; -- 14
        TB : OUT STD_LOGIC; -- 15
        TA : OUT STD_LOGIC; -- 16
        TD : OUT STD_LOGIC; -- 17
        PL : OUT STD_LOGIC; -- 18
        PI : OUT STD_LOGIC; -- 19
        IL : OUT STD_LOGIC; -- 20
        MC : OUT STD_LOGIC; -- 21
        MS : OUT STD_LOGIC_VECTOR(2 DOWNTO 0); -- 22 to 24
        NA : OUT STD_LOGIC_VECTOR(16 DOWNTO 0) -- 25 to 41
    );
END ctrl_mem;

ARCHITECTURE Behavioral OF ctrl_mem IS
    -- we will use the least significant 8 bit of the IN_CAR - array(0 to 255)
    TYPE mem_array IS ARRAY(0 TO 255) OF STD_LOGIC_VECTOR(41 DOWNTO 0);
    -- initialise the control memory
    SIGNAL control_mem : mem_array := (
        -- |41 25|24 22|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
        -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
        -- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
        "000000000000000000000000000000000000000000", -- 0
        "000000000000000010000000000000000000000000", -- 1
        "000000000000000100000000000000000000000000", -- 2
        "000000000000000110000000000000000000000000", -- 3
        "000000000000001000000000000000000000000000", -- 4
        "000000000000001010000000000000000000000000", -- 5
        "000000000000001100000000000000000000000000", -- 6
        "000000000000001110000000000000000000000000", -- 7
        "000000000000010000000000000000000000000000", -- 8
        "000000000000010010000000000000000000000000", -- 9
        "000000000000010100000000000000000000000000", -- a
        "000000000000010110000000000000000000000000", -- b
        "000000000000011000000000000000000000000000", -- c
        "000000000000011010000000000000000000000000", -- d
        "000000000000011100000000000000000000000000", -- e
        "000000000000011110000000000000000000000000", -- f
        "000000000000100000000000000000000000000000", -- 10
        "000000000000100010000000000000000000000000", -- 11
        "000000000000100100000000000000000000000000", -- 12
        "000000000000100110000000000000000000000000", -- 13
        "000000000000101000000000000000000000000000", -- 14
        "000000000000101010000000000000000000000000", -- 15
        "000000000000101100000000000000000000000000", -- 16
        "000000000000101110000000000000000000000000", -- 17
        "000000000000110000000000000000000000000000", -- 18
        "000000000000110010000000000000000000000000", -- 19
        "000000000000110100000000000000000000000000", -- 1a
        "000000000000110110000000000000000000000000", -- 1b
        "000000000000111000000000000000000000000000", -- 1c
        "000000000000111010000000000000000000000000", -- 1d
        "000000000000111100000000000000000000000000", -- 1e
        "000000000000111110000000000000000000000000", -- 1f
        "000000000001000000000000000000000000000000", -- 20
        "000000000001000010000000000000000000000000", -- 21
        "000000000001000100000000000000000000000000", -- 22
        "000000000001000110000000000000000000000000", -- 23
        "000000000001001000000000000000000000000000", -- 24
        "000000000001001010000000000000000000000000", -- 25
        "000000000001001100000000000000000000000000", -- 26
        "000000000001001110000000000000000000000000", -- 27
        "000000000001010000000000000000000000000000", -- 28
        "000000000001010010000000000000000000000000", -- 29
        "000000000001010100000000000000000000000000", -- 2a
        "000000000001010110000000000000000000000000", -- 2b
        "000000000001011000000000000000000000000000", -- 2c
        "000000000001011010000000000000000000000000", -- 2d
        "000000000001011100000000000000000000000000", -- 2e
        "000000000001011110000000000000000000000000", -- 2f
        "000000000001100000000000000000000000000000", -- 30
        "000000000001100010000000000000000000000000", -- 31
        "000000000001100100000000000000000000000000", -- 32
        "000000000001100110000000000000000000000000", -- 33
        "000000000001101000000000000000000000000000", -- 34
        "000000000001101010000000000000000000000000", -- 35
        "000000000001101100000000000000000000000000", -- 36
        "000000000001101110000000000000000000000000", -- 37
        "000000000001110000000000000000000000000000", -- 38
        "000000000001110010000000000000000000000000", -- 39
        "000000000001110100000000000000000000000000", -- 3a
        "000000000001110110000000000000000000000000", -- 3b
        "000000000001111000000000000000000000000000", -- 3c
        "000000000001111010000000000000000000000000", -- 3d
        "000000000001111100000000000000000000000000", -- 3e
        "000000000001111110000000000000000000000000", -- 3f
        "000000000010000000000000000000000000000000", -- 40
        "000000000010000010000000000000000000000000", -- 41
        "000000000010000100000000000000000000000000", -- 42
        "000000000010000110000000000000000000000000", -- 43
        "000000000010001000000000000000000000000000", -- 44
        "000000000010001010000000000000000000000000", -- 45
        "000000000010001100000000000000000000000000", -- 46
        "000000000010001110000000000000000000000000", -- 47
        "000000000010010000000000000000000000000000", -- 48
        "000000000010010010000000000000000000000000", -- 49
        "000000000010010100000000000000000000000000", -- 4a
        "000000000010010110000000000000000000000000", -- 4b
        "000000000010011000000000000000000000000000", -- 4c
        "000000000010011010000000000000000000000000", -- 4d
        "000000000010011100000000000000000000000000", -- 4e
        "000000000010011110000000000000000000000000", -- 4f
        "000000000010100000000000000000000000000000", -- 50
        "000000000010100010000000000000000000000000", -- 51
        "000000000010100100000000000000000000000000", -- 52
        "000000000010100110000000000000000000000000", -- 53
        "000000000010101000000000000000000000000000", -- 54
        "000000000010101010000000000000000000000000", -- 55
        "000000000010101100000000000000000000000000", -- 56
        "000000000010101110000000000000000000000000", -- 57
        "000000000010110000000000000000000000000000", -- 58
        "000000000010110010000000000000000000000000", -- 59
        "000000000010110100000000000000000000000000", -- 5a
        "000000000010110110000000000000000000000000", -- 5b
        "000000000010111000000000000000000000000000", -- 5c
        "000000000010111010000000000000000000000000", -- 5d
        "000000000010111100000000000000000000000000", -- 5e
        "000000000010111110000000000000000000000000", -- 5f
        "000000000011000000000000000000000000000000", -- 60
        "000000000011000010000000000000000000000000", -- 61
        "000000000011000100000000000000000000000000", -- 62
        "000000000011000110000000000000000000000000", -- 63
        "000000000011001000000000000000000000000000", -- 64
        "000000000011001010000000000000000000000000", -- 65
        "000000000011001100000000000000000000000000", -- 66
        "000000000011001110000000000000000000000000", -- 67
        "000000000011010000000000000000000000000000", -- 68
        "000000000011010010000000000000000000000000", -- 69
        "000000000011010100000000000000000000000000", -- 6a
        "000000000011010110000000000000000000000000", -- 6b
        "000000000011011000000000000000000000000000", -- 6c
        "000000000011011010000000000000000000000000", -- 6d
        "000000000011011100000000000000000000000000", -- 6e
        "000000000011011110000000000000000000000000", -- 6f
        "000000000011100000000000000000000000000000", -- 70
        "000000000011100010000000000000000000000000", -- 71
        "000000000011100100000000000000000000000000", -- 72
        "000000000011100110000000000000000000000000", -- 73
        "000000000011101000000000000000000000000000", -- 74
        "000000000011101010000000000000000000000000", -- 75
        "000000000011101100000000000000000000000000", -- 76
        "000000000011101110000000000000000000000000", -- 77
        "000000000011110000000000000000000000000000", -- 78
        "000000000011110010000000000000000000000000", -- 79
        "000000000011110100000000000000000000000000", -- 7a
        "000000000011110110000000000000000000000000", -- 7b
        "000000000011111000000000000000000000000000", -- 7c
        "000000000011111010000000000000000000000000", -- 7d
        "000000000011111100000000000000000000000000", -- 7e
        "000000000011111110000000000000000000000000", -- 7f
        "000000000100000000000000000000000000000000", -- 80
        "000000000100000010000000000000000000000000", -- 81
        "000000000100000100000000000000000000000000", -- 82
        "000000000100000110000000000000000000000000", -- 83
        "000000000100001000000000000000000000000000", -- 84
        "000000000100001010000000000000000000000000", -- 85
        "000000000100001100000000000000000000000000", -- 86
        "000000000100001110000000000000000000000000", -- 87
        "000000000100010000000000000000000000000000", -- 88
        "000000000100010010000000000000000000000000", -- 89
        "000000000100010100000000000000000000000000", -- 8a
        "000000000100010110000000000000000000000000", -- 8b
        "000000000100011000000000000000000000000000", -- 8c
        "000000000100011010000000000000000000000000", -- 8d
        "000000000100011100000000000000000000000000", -- 8e
        "000000000100011110000000000000000000000000", -- 8f
        "000000000100100000000000000000000000000000", -- 90
        "000000000100100010000000000000000000000000", -- 91
        "000000000100100100000000000000000000000000", -- 92
        "000000000100100110000000000000000000000000", -- 93
        "000000000100101000000000000000000000000000", -- 94
        "000000000100101010000000000000000000000000", -- 95
        "000000000100101100000000000000000000000000", -- 96
        "000000000100101110000000000000000000000000", -- 97
        "000000000100110000000000000000000000000000", -- 98
        "000000000100110010000000000000000000000000", -- 99
        "000000000100110100000000000000000000000000", -- 9a
        "000000000100110110000000000000000000000000", -- 9b
        "000000000100111000000000000000000000000000", -- 9c
        "000000000100111010000000000000000000000000", -- 9d
        "000000000100111100000000000000000000000000", -- 9e
        "000000000100111110000000000000000000000000", -- 9f
        "000000000101000000000000000000000000000000", -- a0
        "000000000101000010000000000000000000000000", -- a1
        "000000000101000100000000000000000000000000", -- a2
        "000000000101000110000000000000000000000000", -- a3
        "000000000101001000000000000000000000000000", -- a4
        "000000000101001010000000000000000000000000", -- a5
        "000000000101001100000000000000000000000000", -- a6
        "000000000101001110000000000000000000000000", -- a7
        "000000000101010000000000000000000000000000", -- a8
        "000000000101010010000000000000000000000000", -- a9
        "000000000101010100000000000000000000000000", -- aa
        "000000000101010110000000000000000000000000", -- ab
        "000000000101011000000000000000000000000000", -- ac
        "000000000101011010000000000000000000000000", -- ad
        "000000000101011100000000000000000000000000", -- ae
        "000000000101011110000000000000000000000000", -- af
        "000000000101100000000000000000000000000000", -- b0
        "000000000101100010000000000000000000000000", -- b1
        "000000000101100100000000000000000000000000", -- b2
        "000000000101100110000000000000000000000000", -- b3
        "000000000101101000000000000000000000000000", -- b4
        "000000000101101010000000000000000000000000", -- b5
        "000000000101101100000000000000000000000000", -- b6
        "000000000101101110000000000000000000000000", -- b7
        "000000000101110000000000000000000000000000", -- b8
        "000000000101110010000000000000000000000000", -- b9
        "000000000101110100000000000000000000000000", -- ba
        "000000000101110110000000000000000000000000", -- bb
        "000000000101111000000000000000000000000000", -- bc
        "000000000101111010000000000000000000000000", -- bd
        "000000000101111100000000000000000000000000", -- be
        "000000000101111110000000000000000000000000", -- bf
        "000000000110000000000000000000000000000000", -- c0
        "000000000110000010000000000000000000000000", -- c1
        "000000000110000100000000000000000000000000", -- c2
        "000000000110000110000000000000000000000000", -- c3
        "000000000110001000000000000000000000000000", -- c4
        "000000000110001010000000000000000000000000", -- c5
        "000000000110001100000000000000000000000000", -- c6
        "000000000110001110000000000000000000000000", -- c7
        "000000000110010000000000000000000000000000", -- c8
        "000000000110010010000000000000000000000000", -- c9
        "000000000110010100000000000000000000000000", -- ca
        "000000000110010110000000000000000000000000", -- cb
        "000000000110011000000000000000000000000000", -- cc
        "000000000110011010000000000000000000000000", -- cd
        "000000000110011100000000000000000000000000", -- ce
        "000000000110011110000000000000000000000000", -- cf
        "000000000110100000000000000000000000000000", -- d0
        "000000000110100010000000000000000000000000", -- d1
        "000000000110100100000000000000000000000000", -- d2
        "000000000110100110000000000000000000000000", -- d3
        "000000000110101000000000000000000000000000", -- d4
        "000000000110101010000000000000000000000000", -- d5
        "000000000110101100000000000000000000000000", -- d6
        "000000000110101110000000000000000000000000", -- d7
        "000000000110110000000000000000000000000000", -- d8
        "000000000110110010000000000000000000000000", -- d9
        "000000000110110100000000000000000000000000", -- da
        "000000000110110110000000000000000000000000", -- db
        "000000000110111000000000000000000000000000", -- dc
        "000000000110111010000000000000000000000000", -- dd
        "000000000110111100000000000000000000000000", -- de
        "000000000110111110000000000000000000000000", -- df
        "000000000111000000000000000000000000000000", -- e0
        "000000000111000010000000000000000000000000", -- e1
        "000000000111000100000000000000000000000000", -- e2
        "000000000111000110000000000000000000000000", -- e3
        "000000000111001000000000000000000000000000", -- e4
        "000000000111001010000000000000000000000000", -- e5
        "000000000111001100000000000000000000000000", -- e6
        "000000000111001110000000000000000000000000", -- e7
        "000000000111010000000000000000000000000000", -- e8
        "000000000111010010000000000000000000000000", -- e9
        "000000000111010100000000000000000000000000", -- ea
        "000000000111010110000000000000000000000000", -- eb
        "000000000111011000000000000000000000000000", -- ec
        "000000000111011010000000000000000000000000", -- ed
        "000000000111011100000000000000000000000000", -- ee
        "000000000111011110000000000000000000000000", -- ef
        "000000000111100000000000000000000000000000", -- f0
        "000000000111100010000000000000000000000000", -- f1
        "000000000111100100000000000000000000000000", -- f2
        "000000000111100110000000000000000000000000", -- f3
        "000000000111101000000000000000000000000000", -- f4
        "000000000111101010000000000000000000000000", -- f5
        "000000000111101100000000000000000000000000", -- f6
        "000000000111101110000000000000000000000000", -- f7
        "000000000111110000000000000000000000000000", -- f8
        "000000000111110010000000000000000000000000", -- f9
        "000000000111110100000000000000000000000000", -- fa
        "000000000111110110000000000000000000000000", -- fb
        "000000000111111000000000000000000000000000", -- fc
        "000000000111111010000000000000000000000000", -- fd
        "000000000111111100000000000000000000000000", -- fe
        "000000000111111110000000000000000000000000" -- ff
    );
    SIGNAL adrs_content : STD_LOGIC_VECTOR(41 DOWNTO 0);

BEGIN
    adrs_content <= control_mem(to_integer(unsigned(IN_CAR(8 DOWNTO 0)))) AFTER 2ns;
    FL <= adrs_content(0); -- 0
    RZ <= adrs_content(1); -- 1
    RN <= adrs_content(2); -- 2
    RC <= adrs_content(3); -- 3
    RV <= adrs_content(4); -- 4
    MW <= adrs_content(5); -- 5
    MM <= adrs_content(6); -- 6
    RW <= adrs_content(7); -- 7
    MD <= adrs_content(8); -- 8
    FS <= adrs_content(13 DOWNTO 9); -- 9 to 13
    MB <= adrs_content(14); -- 14
    TB <= adrs_content(15); -- 15
    TA <= adrs_content(16); -- 16
    TD <= adrs_content(17); -- 17
    PL <= adrs_content(18); -- 18
    PI <= adrs_content(19); -- 19
    IL <= adrs_content(20); -- 20
    MC <= adrs_content(21); -- 21
    MS <= adrs_content(24 DOWNTO 22); -- 22 to 24
    NA <= adrs_content(41 DOWNTO 25); -- 25 to 41
END Behavioral;