LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY memory_512 IS
    PORT (
        mem_address : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_in : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        write_enable, clk : IN STD_LOGIC;
        data_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END memory_512;

ARCHITECTURE Behavioral OF memory_512 IS
    TYPE mem_array IS ARRAY(0 TO 511) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL memory_512 : mem_array := (
        x"00000000", x"00000001", x"00000002", x"00000003", x"00000004", x"00000005", x"00000006", x"00000007",
        x"00000008", x"00000009", x"0000000a", x"0000000b", x"0000000c", x"0000000d", x"0000000e", x"0000000f",
        x"00000010", x"00000011", x"00000012", x"00000013", x"00000014", x"00000015", x"00000016", x"00000017",
        x"00000018", x"00000019", x"0000001a", x"0000001b", x"0000001c", x"0000001d", x"0000001e", x"0000001f",
        x"00000020", x"00000021", x"00000022", x"00000023", x"00000024", x"00000025", x"00000026", x"00000027",
        x"00000028", x"00000029", x"0000002a", x"0000002b", x"0000002c", x"0000002d", x"0000002e", x"0000002f",
        x"00000030", x"00000031", x"00000032", x"00000033", x"00000034", x"00000035", x"00000036", x"00000037",
        x"00000038", x"00000039", x"0000003a", x"0000003b", x"0000003c", x"0000003d", x"0000003e", x"0000003f",
        x"00000040", x"00000041", x"00000042", x"00000043", x"00000044", x"00000045", x"00000046", x"00000047",
        x"00000048", x"00000049", x"0000004a", x"0000004b", x"0000004c", x"0000004d", x"0000004e", x"0000004f",
        x"00000050", x"00000051", x"00000052", x"00000053", x"00000054", x"00000055", x"00000056", x"00000057",
        x"00000058", x"00000059", x"0000005a", x"0000005b", x"0000005c", x"0000005d", x"0000005e", x"0000005f",
        x"00000060", x"00000061", x"00000062", x"00000063", x"00000064", x"00000065", x"00000066", x"00000067",
        x"00000068", x"00000069", x"0000006a", x"0000006b", x"0000006c", x"0000006d", x"0000006e", x"0000006f",
        x"00000070", x"00000071", x"00000072", x"00000073", x"00000074", x"00000075", x"00000076", x"00000077",
        x"00000078", x"00000079", x"0000007a", x"0000007b", x"0000007c", x"0000007d", x"0000007e", x"0000007f",
        x"00000080", x"00000081", x"00000082", x"00000083", x"00000084", x"00000085", x"00000086", x"00000087",
        x"00000088", x"00000089", x"0000008a", x"0000008b", x"0000008c", x"0000008d", x"0000008e", x"0000008f",
        x"00000090", x"00000091", x"00000092", x"00000093", x"00000094", x"00000095", x"00000096", x"00000097",
        x"00000098", x"00000099", x"0000009a", x"0000009b", x"0000009c", x"0000009d", x"0000009e", x"0000009f",
        x"000000a0", x"000000a1", x"000000a2", x"000000a3", x"000000a4", x"000000a5", x"000000a6", x"000000a7",
        x"000000a8", x"000000a9", x"000000aa", x"000000ab", x"000000ac", x"000000ad", x"000000ae", x"000000af",
        x"000000b0", x"000000b1", x"000000b2", x"000000b3", x"000000b4", x"000000b5", x"000000b6", x"000000b7",
        x"000000b8", x"000000b9", x"000000ba", x"000000bb", x"000000bc", x"000000bd", x"000000be", x"000000bf",
        x"000000c0", x"000000c1", x"000000c2", x"000000c3", x"000000c4", x"000000c5", x"000000c6", x"000000c7",
        x"000000c8", x"000000c9", x"000000ca", x"000000cb", x"000000cc", x"000000cd", x"000000ce", x"000000cf",
        x"000000d0", x"000000d1", x"000000d2", x"000000d3", x"000000d4", x"000000d5", x"000000d6", x"000000d7",
        x"000000d8", x"000000d9", x"000000da", x"000000db", x"000000dc", x"000000dd", x"000000de", x"000000df",
        x"000000e0", x"000000e1", x"000000e2", x"000000e3", x"000000e4", x"000000e5", x"000000e6", x"000000e7",
        x"000000e8", x"000000e9", x"000000ea", x"000000eb", x"000000ec", x"000000ed", x"000000ee", x"000000ef",
        x"000000f0", x"000000f1", x"000000f2", x"000000f3", x"000000f4", x"000000f5", x"000000f6", x"000000f7",
        x"000000f8", x"000000f9", x"000000fa", x"000000fb", x"000000fc", x"000000fd", x"000000fe", x"000000ff",
        x"00000100", x"00000101", x"00000102", x"00000103", x"00000104", x"00000105", x"00000106", x"00000107",
        x"00000108", x"00000109", x"0000010a", x"0000010b", x"0000010c", x"0000010d", x"0000010e", x"0000010f",
        x"00000110", x"00000111", x"00000112", x"00000113", x"00000114", x"00000115", x"00000116", x"00000117",
        x"00000118", x"00000119", x"0000011a", x"0000011b", x"0000011c", x"0000011d", x"0000011e", x"0000011f",
        x"00000120", x"00000121", x"00000122", x"00000123", x"00000124", x"00000125", x"00000126", x"00000127",
        x"00000128", x"00000129", x"0000012a", x"0000012b", x"0000012c", x"0000012d", x"0000012e", x"0000012f",
        x"00000130", x"00000131", x"00000132", x"00000133", x"00000134", x"00000135", x"00000136", x"00000137",
        x"00000138", x"00000139", x"0000013a", x"0000013b", x"0000013c", x"0000013d", x"0000013e", x"0000013f",
        x"00000140", x"00000141", x"00000142", x"00000143", x"00000144", x"00000145", x"00000146", x"00000147",
        x"00000148", x"00000149", x"0000014a", x"0000014b", x"0000014c", x"0000014d", x"0000014e", x"0000014f",
        x"00000150", x"00000151", x"00000152", x"00000153", x"00000154", x"00000155", x"00000156", x"00000157",
        x"00000158", x"00000159", x"0000015a", x"0000015b", x"0000015c", x"0000015d", x"0000015e", x"0000015f",
        x"00000160", x"00000161", x"00000162", x"00000163", x"00000164", x"00000165", x"00000166", x"00000167",
        x"00000168", x"00000169", x"0000016a", x"0000016b", x"0000016c", x"0000016d", x"0000016e", x"0000016f",
        x"00000170", x"00000171", x"00000172", x"00000173", x"00000174", x"00000175", x"00000176", x"00000177",
        x"00000178", x"00000179", x"0000017a", x"0000017b", x"0000017c", x"0000017d", x"0000017e", x"0000017f",
        x"00000180", x"00000181", x"00000182", x"00000183", x"00000184", x"00000185", x"00000186", x"00000187",
        x"00000188", x"00000189", x"0000018a", x"0000018b", x"0000018c", x"0000018d", x"0000018e", x"0000018f",
        x"00000190", x"00000191", x"00000192", x"00000193", x"00000194", x"00000195", x"00000196", x"00000197",
        x"00000198", x"00000199", x"0000019a", x"0000019b", x"0000019c", x"0000019d", x"0000019e", x"0000019f",
        x"000001a0", x"000001a1", x"000001a2", x"000001a3", x"000001a4", x"000001a5", x"000001a6", x"000001a7",
        x"000001a8", x"000001a9", x"000001aa", x"000001ab", x"000001ac", x"000001ad", x"000001ae", x"000001af",
        x"000001b0", x"000001b1", x"000001b2", x"000001b3", x"000001b4", x"000001b5", x"000001b6", x"000001b7",
        x"000001b8", x"000001b9", x"000001ba", x"000001bb", x"000001bc", x"000001bd", x"000001be", x"000001bf",
        x"000001c0", x"000001c1", x"000001c2", x"000001c3", x"000001c4", x"000001c5", x"000001c6", x"000001c7",
        x"000001c8", x"000001c9", x"000001ca", x"000001cb", x"000001cc", x"000001cd", x"000001ce", x"000001cf",
        x"000001d0", x"000001d1", x"000001d2", x"000001d3", x"000001d4", x"000001d5", x"000001d6", x"000001d7",
        x"000001d8", x"000001d9", x"000001da", x"000001db", x"000001dc", x"000001dd", x"000001de", x"000001df",
        x"000001e0", x"000001e1", x"000001e2", x"000001e3", x"000001e4", x"000001e5", x"000001e6", x"000001e7",
        x"000001e8", x"000001e9", x"000001ea", x"000001eb", x"000001ec", x"000001ed", x"000001ee", x"000001ef",
        x"000001f0", x"000001f1", x"000001f2", x"000001f3", x"000001f4", x"000001f5", x"000001f6", x"000001f7",
        x"000001f8", x"000001f9", x"000001fa", x"000001fb", x"000001fc", x"000001fd", x"000001fe", x"000001ff"
    );

BEGIN
    mem_process : process(clk)
    begin
        if (rising_edge(clk)) then
            if (write_enable = '1') then 
                memory_512(to_integer(unsigned(mem_address(8 DOWNTO 0)))) <= data_in after 1 ns;
            end if;
        end if;
    end process ; -- mem_process
    data_out <= memory_512(to_integer(unsigned(mem_address(8 DOWNTO 0)))) after 1 ns WHEN write_enable = '0';
END Behavioral;