LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux32_tb IS
END mux32_tb;

ARCHITECTURE Behavioral OF mux32_tb IS
    COMPONENT mux32
        PORT (
            in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12,
            in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23,
            in24, in25, in26, in27, in28, in29, in30, in31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            s0, s1, s2, s3, s4 : IN STD_LOGIC;
            z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
        );
    END COMPONENT;

    -- input
    SIGNAL in0 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in1 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in2 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in3 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in4 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in5 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in6 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in7 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in8 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in9 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in10 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in11 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in12 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in13 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in14 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in15 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in16 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in17 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in18 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in19 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in20 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in21 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in22 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in23 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in24 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in25 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in26 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in27 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in28 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in29 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in30 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in31 : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');

    SIGNAL s0 : STD_LOGIC := '0';
    SIGNAL s1 : STD_LOGIC := '0';
    SIGNAL s2 : STD_LOGIC := '0';
    SIGNAL s3 : STD_LOGIC := '0';
    SIGNAL s4 : STD_LOGIC := '0';

    -- output
    SIGNAL Z : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
BEGIN
    uut : mux32 PORT MAP(
        in0 => in0, in1 => in1, in2 => in2, in3 => in3, in4 => in4, in5 => in5, in6 => in6, in7 => in7, in8 => in8, in9 => in9, in10 => in10, in11 => in11,
        in12 => in12, in13 => in13, in14 => in14, in15 => in15, in16 => in16, in17 => in17, in18 => in18, in19 => in19, in20 => in20, in21 => in21, in22 => in22,
        in23 => in23, in24 => in24, in25 => in25, in26 => in26, in27 => in27, in28 => in28, in29 => in29, in30 => in30, in31 => in31,
        s0 => s0, s1 => s1, s2 => s2, s3 => s3, s4 => s4,
        Z => Z
    );
    stim_proc : PROCESS
    BEGIN
        in0 <= "00000000000000000000000000000111";
        in1 <= "00000000000000000000000000001110";
        in2 <= "00000000000000000000000000011100";
        in3 <= "00000000000000000000000000111000";
        in4 <= "00000000000000000000000001110000";
        in5 <= "00000000000000000000000011100000";
        in6 <= "00000000000000000000000111000000";
        in7 <= "00000000000000000000001110000000";
        in8 <= "00000000000000000000011100000000";
        in9 <= "00000000000000000000111000000000";
        in10 <= "00000000000000000001110000000000";
        in11 <= "00000000000000000011100000000000";
        in12 <= "00000000000000000111000000000000";
        in13 <= "00000000000000001110000000000000";
        in14 <= "00000000000000011100000000000000";
        in15 <= "00000000000000111000000000000000";
        in16 <= "00000000000001110000000000000000";
        in17 <= "00000000000011100000000000000000";
        in18 <= "00000000000111000000000000000000";
        in19 <= "00000000001110000000000000000000";
        in20 <= "00000000011100000000000000000000";
        in21 <= "00000000111000000000000000000000";
        in22 <= "00000001110000000000000000000000";
        in23 <= "00000011100000000000000000000000";
        in24 <= "00000111000000000000000000000000";
        in25 <= "00001110000000000000000000000000";
        in26 <= "00011100000000000000000000000000";
        in27 <= "00111000000000000000000000000000";
        in28 <= "01110000000000000000000000000000";
        in29 <= "11100000000000000000000000000000";
        in30 <= "11000000000000000000000000000000";
        in31 <= "10000000000000000000000000000000";

        s0 <= '0';
        s1 <= '0';
        s2 <= '0';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '0';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '0';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '0';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '1';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '1';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '1';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '0';
        s2 <= '1';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '0';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '0';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '0';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '0';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '1';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '1';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '1';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '0';
        s1 <= '1';
        s2 <= '1';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '0';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '0';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '0';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '0';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '1';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '1';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '1';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '0';
        s2 <= '1';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '0';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '0';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '0';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '0';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '1';
        s3 <= '0';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '1';
        s3 <= '0';
        s4 <= '1';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '1';
        s3 <= '1';
        s4 <= '0';
        WAIT FOR 5ns;
        s0 <= '1';
        s1 <= '1';
        s2 <= '1';
        s3 <= '1';
        s4 <= '1';
        WAIT FOR 5ns;
    END PROCESS;
END Behavioral;